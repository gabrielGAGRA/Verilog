module porta_e(
    input a,
    input b,
    output y
);
    assign y = a & b;
endmodule
